module ALU(
  input         clock,
  input         reset,
  input  [31:0] io_op1,
  input  [31:0] io_op2,
  input  [3:0]  io_sel,
  output [31:0] io_result,
  output        io_cmpResult
);
  wire  _T = 4'h0 == io_sel; // @[Conditional.scala 37:30]
  wire [31:0] _T_2 = io_op1 + io_op2; // @[ALU.scala 19:36]
  wire  _T_3 = 4'h1 == io_sel; // @[Conditional.scala 37:30]
  wire [31:0] _T_5 = io_op1 - io_op2; // @[ALU.scala 20:36]
  wire  _T_6 = 4'h2 == io_sel; // @[Conditional.scala 37:30]
  wire [63:0] _T_7 = io_op1 * io_op2; // @[ALU.scala 21:36]
  wire  _T_8 = 4'h3 == io_sel; // @[Conditional.scala 37:30]
  wire [31:0] _T_10 = io_op1 + 32'h1; // @[ALU.scala 22:36]
  wire  _T_11 = 4'h4 == io_sel; // @[Conditional.scala 37:30]
  wire [31:0] _T_13 = io_op1 - 32'h1; // @[ALU.scala 23:36]
  wire  _T_14 = 4'h5 == io_sel; // @[Conditional.scala 37:30]
  wire [31:0] _T_15 = ~io_op1; // @[ALU.scala 24:29]
  wire  _T_16 = 4'h6 == io_sel; // @[Conditional.scala 37:30]
  wire [31:0] _T_17 = io_op1 & io_op2; // @[ALU.scala 25:36]
  wire  _T_18 = 4'h7 == io_sel; // @[Conditional.scala 37:30]
  wire [31:0] _T_19 = io_op1 | io_op2; // @[ALU.scala 26:36]
  wire  _T_20 = 4'h8 == io_sel; // @[Conditional.scala 37:30]
  wire [31:0] _T_21 = io_op1 ^ io_op2; // @[ALU.scala 27:36]
  wire  _T_22 = 4'h9 == io_sel; // @[Conditional.scala 37:30]
  wire  _T_23 = io_op1 == io_op2; // @[ALU.scala 30:39]
  wire  _T_24 = 4'ha == io_sel; // @[Conditional.scala 37:30]
  wire  _T_25 = io_op1 != io_op2; // @[ALU.scala 31:40]
  wire  _T_26 = 4'hb == io_sel; // @[Conditional.scala 37:30]
  wire  _T_27 = io_op1 > io_op2; // @[ALU.scala 32:40]
  wire  _T_28 = 4'hc == io_sel; // @[Conditional.scala 37:30]
  wire  _T_29 = io_op1 >= io_op2; // @[ALU.scala 33:40]
  wire  _T_30 = 4'hd == io_sel; // @[Conditional.scala 37:30]
  wire  _T_31 = io_op1 < io_op2; // @[ALU.scala 34:40]
  wire  _T_32 = 4'he == io_sel; // @[Conditional.scala 37:30]
  wire  _T_33 = io_op1 <= io_op2; // @[ALU.scala 35:40]
  wire  _T_34 = 4'hf == io_sel; // @[Conditional.scala 37:30]
  wire  _GEN_1 = _T_32 ? _T_33 : _T_34; // @[Conditional.scala 39:67]
  wire  _GEN_2 = _T_30 ? _T_31 : _GEN_1; // @[Conditional.scala 39:67]
  wire  _GEN_3 = _T_28 ? _T_29 : _GEN_2; // @[Conditional.scala 39:67]
  wire  _GEN_4 = _T_26 ? _T_27 : _GEN_3; // @[Conditional.scala 39:67]
  wire  _GEN_5 = _T_24 ? _T_25 : _GEN_4; // @[Conditional.scala 39:67]
  wire  _GEN_6 = _T_22 ? _T_23 : _GEN_5; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_7 = _T_20 ? _T_21 : 32'h0; // @[Conditional.scala 39:67]
  wire  _GEN_8 = _T_20 ? 1'h0 : _GEN_6; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_9 = _T_18 ? _T_19 : _GEN_7; // @[Conditional.scala 39:67]
  wire  _GEN_10 = _T_18 ? 1'h0 : _GEN_8; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_11 = _T_16 ? _T_17 : _GEN_9; // @[Conditional.scala 39:67]
  wire  _GEN_12 = _T_16 ? 1'h0 : _GEN_10; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_13 = _T_14 ? _T_15 : _GEN_11; // @[Conditional.scala 39:67]
  wire  _GEN_14 = _T_14 ? 1'h0 : _GEN_12; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_15 = _T_11 ? _T_13 : _GEN_13; // @[Conditional.scala 39:67]
  wire  _GEN_16 = _T_11 ? 1'h0 : _GEN_14; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_17 = _T_8 ? _T_10 : _GEN_15; // @[Conditional.scala 39:67]
  wire  _GEN_18 = _T_8 ? 1'h0 : _GEN_16; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_19 = _T_6 ? _T_7 : {{32'd0}, _GEN_17}; // @[Conditional.scala 39:67]
  wire  _GEN_20 = _T_6 ? 1'h0 : _GEN_18; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_21 = _T_3 ? {{32'd0}, _T_5} : _GEN_19; // @[Conditional.scala 39:67]
  wire  _GEN_22 = _T_3 ? 1'h0 : _GEN_20; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_23 = _T ? {{32'd0}, _T_2} : _GEN_21; // @[Conditional.scala 40:58]
  assign io_result = _GEN_23[31:0]; // @[ALU.scala 14:13 ALU.scala 19:26 ALU.scala 20:26 ALU.scala 21:26 ALU.scala 22:26 ALU.scala 23:26 ALU.scala 24:26 ALU.scala 25:26 ALU.scala 26:26 ALU.scala 27:26]
  assign io_cmpResult = _T ? 1'h0 : _GEN_22; // @[ALU.scala 15:16 ALU.scala 30:29 ALU.scala 31:30 ALU.scala 32:30 ALU.scala 33:30 ALU.scala 34:30 ALU.scala 35:30 ALU.scala 36:30]
endmodule
